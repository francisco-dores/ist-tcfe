.OP
R1 1 2 1.02597459645k
R2 3 2 2.02178008702k
R3 2 5 3.03144887426k
R4 5 0 4.13109833342k
R5 5 6 3.09601431108k
R6 0 4 2.01920057699k
R7 7 8  1.02918842978k
Vs 1 0 0.0 ac 1.0 sin(0 1 1k)
Vo 4 7 0
C 6 8 1.01181492800u
Hvd 5 8 Vo 8.09196032190k
Gib 6 3 2 5 7.28538907285m
.ic v(6)=8.61856072253 v(8)=0.000000e+00
.END
